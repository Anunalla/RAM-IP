`ifndef RAM_PARAMS_SVH
`define RAM_PARAMS_SVH

`define ADDR_WIDTH 3
`define DATA_WIDTH 8
`define RAM_SIZE 8

`endif